package RandomPkg is
end RandomPkg ;